library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.display_types.all;

entity SYNC is
port(
	clk : in std_logic;
	gameStarted : in std_logic;
	player1won : in std_logic;
	player2won : in std_logic;
	hsync, vsync :out std_logic;
	r,g,b : out std_logic_vector(3 downto 0);
	player1 : in coordinate_array (0 to MAX_ELEMENTS - 1, 0 to 1);
	player2 : in coordinate_array (0 to MAX_ELEMENTS - 1, 0 to 1);
	apple_position : in coordinate;
	special_position : in coordinate
);
end entity;

architecture main of SYNC is

constant H_SIZE : integer := 1280;
constant H_FP : integer := 48;
constant H_BP : integer := 248;
constant H_SYNCP : integer := 112;
constant H_OFFSET : integer := H_FP + H_BP + H_SYNCP;

constant V_SIZE : integer := 1024;
constant V_FP : integer := 1;
constant V_BP : integer := 38;
constant V_SYNCP : integer := 3;
constant V_OFFSET : integer := V_FP + V_BP + V_SYNCP;


constant BLACK : integer := 0;
constant WHITE : integer := 1;
constant BLUE : integer := 2;
constant RED : integer := 3;
constant GREEN : integer := 66;


signal hpos : integer range 0 to (H_SIZE + H_OFFSET) := 0;
signal vpos : integer range 0 to (V_SIZE + V_OFFSET) := 0;

signal singleAct : std_logic := '1';

constant circleImage : logic_image(0 to 15, 0 to 15) := (('1','1','1','1','1','1','1','1','1','1','1','1','1','1','1','1')
,('1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1')
,('1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1')
,('1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1')
,('1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1')
,('1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1')
,('1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0')
,('1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0')
,('1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0')
,('1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0')
,('1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0')
,('1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1')
,('1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','1')
,('1','1','1','0','0','0','0','0','0','0','0','0','0','0','1','1')
,('1','1','1','1','0','0','0','0','0','0','0','0','0','1','1','1')
,('1','1','1','1','1','1','0','0','0','0','0','1','1','1','1','1'));

constant gameStartImage : coordinate_array (0 to FIXED_SCREEN_ELEMENTS - 1, 0 to 1) := (0 => (6, 18),1 => (7, 18),2 => (8, 18),3 => (9, 18),4 => (10, 18),5 => (11, 18),6 => (12, 18),7 => (13, 18),8 => (14, 18),9 => (15, 18),10 => (16, 18),11 => (17, 18),12 => (18, 18),13 => (20, 18),14 => (21, 18),15 => (31, 18),16 => (32, 18),17 => (34, 18),18 => (35, 18),19 => (36, 18),20 => (37, 18),21 => (38, 18),22 => (39, 18),23 => (40, 18),24 => (41, 18),25 => (42, 18),26 => (43, 18),27 => (44, 18),28 => (45, 18),29 => (46, 18),30 => (48, 18),31 => (49, 18),32 => (59, 18),33 => (60, 18),34 => (62, 18),35 => (63, 18),36 => (64, 18),37 => (65, 18),38 => (66, 18),39 => (67, 18),40 => (68, 18),41 => (69, 18),42 => (70, 18),43 => (71, 18),44 => (72, 18),45 => (73, 18),46 => (74, 18),47 => (6, 19),48 => (7, 19),49 => (8, 19),50 => (9, 19),51 => (10, 19),52 => (11, 19),53 => (12, 19),54 => (13, 19),55 => (14, 19),56 => (15, 19),57 => (16, 19),58 => (17, 19),59 => (18, 19),60 => (20, 19),61 => (21, 19),62 => (22, 19),63 => (31, 19),64 => (32, 19),65 => (34, 19),66 => (35, 19),67 => (36, 19),68 => (37, 19),69 => (38, 19),70 => (39, 19),71 => (40, 19),72 => (41, 19),73 => (42, 19),74 => (43, 19),75 => (44, 19),76 => (45, 19),77 => (46, 19),78 => (48, 19),79 => (49, 19),80 => (57, 19),81 => (58, 19),82 => (59, 19),83 => (60, 19),84 => (62, 19),85 => (63, 19),86 => (64, 19),87 => (65, 19),88 => (66, 19),89 => (67, 19),90 => (68, 19),91 => (69, 19),92 => (70, 19),93 => (71, 19),94 => (72, 19),95 => (73, 19),96 => (74, 19),97 => (6, 20),98 => (7, 20),99 => (20, 20),100 => (21, 20),101 => (22, 20),102 => (23, 20),103 => (31, 20),104 => (32, 20),105 => (34, 20),106 => (35, 20),107 => (45, 20),108 => (46, 20),109 => (48, 20),110 => (49, 20),111 => (56, 20),112 => (57, 20),113 => (58, 20),114 => (59, 20),115 => (62, 20),116 => (63, 20),117 => (6, 21),118 => (7, 21),119 => (20, 21),120 => (21, 21),121 => (22, 21),122 => (23, 21),123 => (24, 21),124 => (31, 21),125 => (32, 21),126 => (34, 21),127 => (35, 21),128 => (45, 21),129 => (46, 21),130 => (48, 21),131 => (49, 21),132 => (54, 21),133 => (55, 21),134 => (56, 21),135 => (57, 21),136 => (62, 21),137 => (63, 21),138 => (6, 22),139 => (7, 22),140 => (20, 22),141 => (21, 22),142 => (23, 22),143 => (24, 22),144 => (25, 22),145 => (31, 22),146 => (32, 22),147 => (34, 22),148 => (35, 22),149 => (45, 22),150 => (46, 22),151 => (48, 22),152 => (49, 22),153 => (52, 22),154 => (53, 22),155 => (54, 22),156 => (55, 22),157 => (56, 22),158 => (62, 22),159 => (63, 22),160 => (6, 23),161 => (7, 23),162 => (20, 23),163 => (21, 23),164 => (24, 23),165 => (25, 23),166 => (26, 23),167 => (31, 23),168 => (32, 23),169 => (34, 23),170 => (35, 23),171 => (45, 23),172 => (46, 23),173 => (48, 23),174 => (49, 23),175 => (51, 23),176 => (52, 23),177 => (53, 23),178 => (54, 23),179 => (62, 23),180 => (63, 23),181 => (64, 23),182 => (65, 23),183 => (66, 23),184 => (67, 23),185 => (68, 23),186 => (69, 23),187 => (70, 23),188 => (71, 23),189 => (72, 23),190 => (73, 23),191 => (74, 23),192 => (6, 24),193 => (7, 24),194 => (8, 24),195 => (9, 24),196 => (10, 24),197 => (11, 24),198 => (12, 24),199 => (13, 24),200 => (14, 24),201 => (15, 24),202 => (16, 24),203 => (17, 24),204 => (18, 24),205 => (20, 24),206 => (21, 24),207 => (25, 24),208 => (26, 24),209 => (27, 24),210 => (31, 24),211 => (32, 24),212 => (34, 24),213 => (35, 24),214 => (36, 24),215 => (37, 24),216 => (38, 24),217 => (39, 24),218 => (40, 24),219 => (41, 24),220 => (42, 24),221 => (43, 24),222 => (44, 24),223 => (45, 24),224 => (46, 24),225 => (48, 24),226 => (49, 24),227 => (50, 24),228 => (51, 24),229 => (52, 24),230 => (53, 24),231 => (62, 24),232 => (63, 24),233 => (64, 24),234 => (65, 24),235 => (66, 24),236 => (67, 24),237 => (68, 24),238 => (69, 24),239 => (70, 24),240 => (71, 24),241 => (72, 24),242 => (73, 24),243 => (74, 24),244 => (6, 25),245 => (7, 25),246 => (8, 25),247 => (9, 25),248 => (10, 25),249 => (11, 25),250 => (12, 25),251 => (13, 25),252 => (14, 25),253 => (15, 25),254 => (16, 25),255 => (17, 25),256 => (18, 25),257 => (20, 25),258 => (21, 25),259 => (26, 25),260 => (27, 25),261 => (28, 25),262 => (31, 25),263 => (32, 25),264 => (34, 25),265 => (35, 25),266 => (36, 25),267 => (37, 25),268 => (38, 25),269 => (39, 25),270 => (40, 25),271 => (41, 25),272 => (42, 25),273 => (43, 25),274 => (44, 25),275 => (45, 25),276 => (46, 25),277 => (48, 25),278 => (49, 25),279 => (50, 25),280 => (51, 25),281 => (52, 25),282 => (53, 25),283 => (54, 25),284 => (55, 25),285 => (62, 25),286 => (63, 25),287 => (17, 26),288 => (18, 26),289 => (20, 26),290 => (21, 26),291 => (27, 26),292 => (28, 26),293 => (29, 26),294 => (31, 26),295 => (32, 26),296 => (34, 26),297 => (35, 26),298 => (45, 26),299 => (46, 26),300 => (48, 26),301 => (49, 26),302 => (53, 26),303 => (54, 26),304 => (55, 26),305 => (56, 26),306 => (62, 26),307 => (63, 26),308 => (17, 27),309 => (18, 27),310 => (20, 27),311 => (21, 27),312 => (28, 27),313 => (29, 27),314 => (30, 27),315 => (31, 27),316 => (32, 27),317 => (34, 27),318 => (35, 27),319 => (45, 27),320 => (46, 27),321 => (48, 27),322 => (49, 27),323 => (55, 27),324 => (56, 27),325 => (57, 27),326 => (62, 27),327 => (63, 27),328 => (17, 28),329 => (18, 28),330 => (20, 28),331 => (21, 28),332 => (29, 28),333 => (30, 28),334 => (31, 28),335 => (32, 28),336 => (34, 28),337 => (35, 28),338 => (45, 28),339 => (46, 28),340 => (48, 28),341 => (49, 28),342 => (56, 28),343 => (57, 28),344 => (58, 28),345 => (59, 28),346 => (62, 28),347 => (63, 28),348 => (6, 29),349 => (7, 29),350 => (8, 29),351 => (9, 29),352 => (10, 29),353 => (11, 29),354 => (12, 29),355 => (13, 29),356 => (14, 29),357 => (15, 29),358 => (16, 29),359 => (17, 29),360 => (18, 29),361 => (20, 29),362 => (21, 29),363 => (30, 29),364 => (31, 29),365 => (32, 29),366 => (34, 29),367 => (35, 29),368 => (45, 29),369 => (46, 29),370 => (48, 29),371 => (49, 29),372 => (57, 29),373 => (58, 29),374 => (59, 29),375 => (60, 29),376 => (62, 29),377 => (63, 29),378 => (64, 29),379 => (65, 29),380 => (66, 29),381 => (67, 29),382 => (68, 29),383 => (69, 29),384 => (70, 29),385 => (71, 29),386 => (72, 29),387 => (73, 29),388 => (74, 29),389 => (6, 30),390 => (7, 30),391 => (8, 30),392 => (9, 30),393 => (10, 30),394 => (11, 30),395 => (12, 30),396 => (13, 30),397 => (14, 30),398 => (15, 30),399 => (16, 30),400 => (17, 30),401 => (18, 30),402 => (20, 30),403 => (21, 30),404 => (31, 30),405 => (32, 30),406 => (34, 30),407 => (35, 30),408 => (45, 30),409 => (46, 30),410 => (48, 30),411 => (49, 30),412 => (59, 30),413 => (60, 30),414 => (62, 30),415 => (63, 30),416 => (64, 30),417 => (65, 30),418 => (66, 30),419 => (67, 30),420 => (68, 30),421 => (69, 30),422 => (70, 30),423 => (71, 30),424 => (72, 30),425 => (73, 30),426 => (74, 30),427 => (16, 34),428 => (17, 34),429 => (18, 34),430 => (20, 34),431 => (21, 34),432 => (22, 34),433 => (24, 34),434 => (25, 34),435 => (26, 34),436 => (28, 34),437 => (29, 34),438 => (30, 34),439 => (32, 34),440 => (34, 34),441 => (35, 34),442 => (36, 34),443 => (38, 34),444 => (40, 34),445 => (42, 34),446 => (43, 34),447 => (44, 34),448 => (47, 34),449 => (48, 34),450 => (49, 34),451 => (51, 34),452 => (52, 34),453 => (53, 34),454 => (55, 34),455 => (56, 34),456 => (57, 34),457 => (59, 34),458 => (60, 34),459 => (61, 34),460 => (63, 34),461 => (64, 34),462 => (65, 34),463 => (16, 35),464 => (18, 35),465 => (20, 35),466 => (22, 35),467 => (24, 35),468 => (28, 35),469 => (32, 35),470 => (34, 35),471 => (36, 35),472 => (38, 35),473 => (39, 35),474 => (40, 35),475 => (42, 35),476 => (47, 35),477 => (52, 35),478 => (55, 35),479 => (57, 35),480 => (59, 35),481 => (61, 35),482 => (64, 35),483 => (16, 36),484 => (17, 36),485 => (20, 36),486 => (21, 36),487 => (24, 36),488 => (25, 36),489 => (28, 36),490 => (29, 36),491 => (30, 36),492 => (32, 36),493 => (34, 36),494 => (36, 36),495 => (38, 36),496 => (39, 36),497 => (40, 36),498 => (42, 36),499 => (43, 36),500 => (47, 36),501 => (48, 36),502 => (49, 36),503 => (52, 36),504 => (55, 36),505 => (56, 36),506 => (57, 36),507 => (59, 36),508 => (60, 36),509 => (64, 36),510 => (16, 37),511 => (20, 37),512 => (22, 37),513 => (24, 37),514 => (30, 37),515 => (32, 37),516 => (34, 37),517 => (36, 37),518 => (38, 37),519 => (40, 37),520 => (42, 37),521 => (49, 37),522 => (52, 37),523 => (55, 37),524 => (57, 37),525 => (59, 37),526 => (61, 37),527 => (64, 37),528 => (16, 38),529 => (20, 38),530 => (22, 38),531 => (24, 38),532 => (25, 38),533 => (26, 38),534 => (28, 38),535 => (29, 38),536 => (30, 38),537 => (32, 38),538 => (34, 38),539 => (35, 38),540 => (36, 38),541 => (38, 38),542 => (40, 38),543 => (42, 38),544 => (43, 38),545 => (44, 38),546 => (47, 38),547 => (48, 38),548 => (49, 38),549 => (52, 38),550 => (55, 38),551 => (57, 38),552 => (59, 38),553 => (61, 38),554 => (64, 38), others => (-1,-1));
constant player1WinsImage : coordinate_array (0 to FIXED_SCREEN_ELEMENTS - 1, 0 to 1) := (0 => (3, 19),1 => (4, 19),2 => (5, 19),3 => (6, 19),4 => (7, 19),5 => (8, 19),6 => (9, 19),7 => (10, 19),8 => (11, 19),9 => (12, 19),10 => (14, 19),11 => (15, 19),12 => (25, 19),13 => (26, 19),14 => (27, 19),15 => (28, 19),16 => (29, 19),17 => (30, 19),18 => (31, 19),19 => (32, 19),20 => (33, 19),21 => (34, 19),22 => (36, 19),23 => (37, 19),24 => (44, 19),25 => (45, 19),26 => (47, 19),27 => (48, 19),28 => (49, 19),29 => (50, 19),30 => (51, 19),31 => (52, 19),32 => (53, 19),33 => (54, 19),34 => (55, 19),35 => (56, 19),36 => (58, 19),37 => (59, 19),38 => (60, 19),39 => (61, 19),40 => (62, 19),41 => (63, 19),42 => (64, 19),43 => (65, 19),44 => (66, 19),45 => (67, 19),46 => (73, 19),47 => (74, 19),48 => (3, 20),49 => (4, 20),50 => (5, 20),51 => (6, 20),52 => (7, 20),53 => (8, 20),54 => (9, 20),55 => (10, 20),56 => (11, 20),57 => (12, 20),58 => (14, 20),59 => (15, 20),60 => (25, 20),61 => (26, 20),62 => (27, 20),63 => (28, 20),64 => (29, 20),65 => (30, 20),66 => (31, 20),67 => (32, 20),68 => (33, 20),69 => (34, 20),70 => (36, 20),71 => (37, 20),72 => (38, 20),73 => (43, 20),74 => (44, 20),75 => (45, 20),76 => (47, 20),77 => (48, 20),78 => (49, 20),79 => (50, 20),80 => (51, 20),81 => (52, 20),82 => (53, 20),83 => (54, 20),84 => (55, 20),85 => (56, 20),86 => (58, 20),87 => (59, 20),88 => (60, 20),89 => (61, 20),90 => (62, 20),91 => (63, 20),92 => (64, 20),93 => (65, 20),94 => (66, 20),95 => (67, 20),96 => (72, 20),97 => (73, 20),98 => (74, 20),99 => (3, 21),100 => (4, 21),101 => (11, 21),102 => (12, 21),103 => (14, 21),104 => (15, 21),105 => (25, 21),106 => (26, 21),107 => (33, 21),108 => (34, 21),109 => (37, 21),110 => (38, 21),111 => (39, 21),112 => (42, 21),113 => (43, 21),114 => (44, 21),115 => (47, 21),116 => (48, 21),117 => (58, 21),118 => (59, 21),119 => (66, 21),120 => (67, 21),121 => (71, 21),122 => (72, 21),123 => (73, 21),124 => (74, 21),125 => (3, 22),126 => (4, 22),127 => (11, 22),128 => (12, 22),129 => (14, 22),130 => (15, 22),131 => (25, 22),132 => (26, 22),133 => (33, 22),134 => (34, 22),135 => (38, 22),136 => (39, 22),137 => (40, 22),138 => (41, 22),139 => (42, 22),140 => (43, 22),141 => (47, 22),142 => (48, 22),143 => (58, 22),144 => (59, 22),145 => (66, 22),146 => (67, 22),147 => (70, 22),148 => (71, 22),149 => (72, 22),150 => (73, 22),151 => (74, 22),152 => (3, 23),153 => (4, 23),154 => (5, 23),155 => (6, 23),156 => (7, 23),157 => (8, 23),158 => (9, 23),159 => (10, 23),160 => (11, 23),161 => (12, 23),162 => (14, 23),163 => (15, 23),164 => (25, 23),165 => (26, 23),166 => (33, 23),167 => (34, 23),168 => (39, 23),169 => (40, 23),170 => (41, 23),171 => (42, 23),172 => (47, 23),173 => (48, 23),174 => (49, 23),175 => (50, 23),176 => (51, 23),177 => (52, 23),178 => (58, 23),179 => (59, 23),180 => (60, 23),181 => (61, 23),182 => (62, 23),183 => (63, 23),184 => (64, 23),185 => (65, 23),186 => (66, 23),187 => (67, 23),188 => (70, 23),189 => (71, 23),190 => (73, 23),191 => (74, 23),192 => (3, 24),193 => (4, 24),194 => (5, 24),195 => (6, 24),196 => (7, 24),197 => (8, 24),198 => (9, 24),199 => (10, 24),200 => (11, 24),201 => (12, 24),202 => (14, 24),203 => (15, 24),204 => (25, 24),205 => (26, 24),206 => (27, 24),207 => (28, 24),208 => (29, 24),209 => (30, 24),210 => (31, 24),211 => (32, 24),212 => (33, 24),213 => (34, 24),214 => (40, 24),215 => (41, 24),216 => (47, 24),217 => (48, 24),218 => (49, 24),219 => (50, 24),220 => (51, 24),221 => (52, 24),222 => (58, 24),223 => (59, 24),224 => (60, 24),225 => (61, 24),226 => (62, 24),227 => (63, 24),228 => (64, 24),229 => (65, 24),230 => (66, 24),231 => (73, 24),232 => (74, 24),233 => (3, 25),234 => (4, 25),235 => (14, 25),236 => (15, 25),237 => (25, 25),238 => (26, 25),239 => (27, 25),240 => (28, 25),241 => (29, 25),242 => (30, 25),243 => (31, 25),244 => (32, 25),245 => (33, 25),246 => (34, 25),247 => (40, 25),248 => (41, 25),249 => (47, 25),250 => (48, 25),251 => (58, 25),252 => (59, 25),253 => (63, 25),254 => (64, 25),255 => (65, 25),256 => (73, 25),257 => (74, 25),258 => (3, 26),259 => (4, 26),260 => (14, 26),261 => (15, 26),262 => (25, 26),263 => (26, 26),264 => (33, 26),265 => (34, 26),266 => (40, 26),267 => (41, 26),268 => (47, 26),269 => (48, 26),270 => (58, 26),271 => (59, 26),272 => (64, 26),273 => (65, 26),274 => (66, 26),275 => (73, 26),276 => (74, 26),277 => (3, 27),278 => (4, 27),279 => (14, 27),280 => (15, 27),281 => (16, 27),282 => (17, 27),283 => (18, 27),284 => (19, 27),285 => (20, 27),286 => (21, 27),287 => (22, 27),288 => (25, 27),289 => (26, 27),290 => (33, 27),291 => (34, 27),292 => (40, 27),293 => (41, 27),294 => (47, 27),295 => (48, 27),296 => (49, 27),297 => (50, 27),298 => (51, 27),299 => (52, 27),300 => (53, 27),301 => (54, 27),302 => (55, 27),303 => (56, 27),304 => (58, 27),305 => (59, 27),306 => (65, 27),307 => (66, 27),308 => (67, 27),309 => (70, 27),310 => (71, 27),311 => (72, 27),312 => (73, 27),313 => (74, 27),314 => (75, 27),315 => (76, 27),316 => (77, 27),317 => (3, 28),318 => (4, 28),319 => (14, 28),320 => (15, 28),321 => (16, 28),322 => (17, 28),323 => (18, 28),324 => (19, 28),325 => (20, 28),326 => (21, 28),327 => (22, 28),328 => (25, 28),329 => (26, 28),330 => (33, 28),331 => (34, 28),332 => (40, 28),333 => (41, 28),334 => (47, 28),335 => (48, 28),336 => (49, 28),337 => (50, 28),338 => (51, 28),339 => (52, 28),340 => (53, 28),341 => (54, 28),342 => (55, 28),343 => (56, 28),344 => (58, 28),345 => (59, 28),346 => (66, 28),347 => (67, 28),348 => (70, 28),349 => (71, 28),350 => (72, 28),351 => (73, 28),352 => (74, 28),353 => (75, 28),354 => (76, 28),355 => (77, 28),356 => (19, 31),357 => (20, 31),358 => (27, 31),359 => (28, 31),360 => (31, 31),361 => (32, 31),362 => (33, 31),363 => (34, 31),364 => (35, 31),365 => (36, 31),366 => (37, 31),367 => (38, 31),368 => (41, 31),369 => (42, 31),370 => (49, 31),371 => (50, 31),372 => (52, 31),373 => (53, 31),374 => (54, 31),375 => (55, 31),376 => (56, 31),377 => (57, 31),378 => (58, 31),379 => (59, 31),380 => (60, 31),381 => (61, 31),382 => (19, 32),383 => (20, 32),384 => (27, 32),385 => (28, 32),386 => (31, 32),387 => (32, 32),388 => (33, 32),389 => (34, 32),390 => (35, 32),391 => (36, 32),392 => (37, 32),393 => (38, 32),394 => (41, 32),395 => (42, 32),396 => (43, 32),397 => (49, 32),398 => (50, 32),399 => (52, 32),400 => (53, 32),401 => (54, 32),402 => (55, 32),403 => (56, 32),404 => (57, 32),405 => (58, 32),406 => (59, 32),407 => (60, 32),408 => (61, 32),409 => (19, 33),410 => (20, 33),411 => (27, 33),412 => (28, 33),413 => (34, 33),414 => (35, 33),415 => (41, 33),416 => (42, 33),417 => (43, 33),418 => (44, 33),419 => (49, 33),420 => (50, 33),421 => (52, 33),422 => (53, 33),423 => (19, 34),424 => (20, 34),425 => (21, 34),426 => (23, 34),427 => (24, 34),428 => (26, 34),429 => (27, 34),430 => (28, 34),431 => (34, 34),432 => (35, 34),433 => (41, 34),434 => (42, 34),435 => (43, 34),436 => (44, 34),437 => (45, 34),438 => (49, 34),439 => (50, 34),440 => (52, 34),441 => (53, 34),442 => (20, 35),443 => (21, 35),444 => (23, 35),445 => (24, 35),446 => (26, 35),447 => (27, 35),448 => (34, 35),449 => (35, 35),450 => (41, 35),451 => (42, 35),452 => (44, 35),453 => (45, 35),454 => (46, 35),455 => (49, 35),456 => (50, 35),457 => (52, 35),458 => (53, 35),459 => (54, 35),460 => (55, 35),461 => (56, 35),462 => (57, 35),463 => (58, 35),464 => (59, 35),465 => (60, 35),466 => (61, 35),467 => (20, 36),468 => (21, 36),469 => (22, 36),470 => (23, 36),471 => (24, 36),472 => (25, 36),473 => (26, 36),474 => (27, 36),475 => (34, 36),476 => (35, 36),477 => (41, 36),478 => (42, 36),479 => (45, 36),480 => (46, 36),481 => (47, 36),482 => (49, 36),483 => (50, 36),484 => (52, 36),485 => (53, 36),486 => (54, 36),487 => (55, 36),488 => (56, 36),489 => (57, 36),490 => (58, 36),491 => (59, 36),492 => (60, 36),493 => (61, 36),494 => (20, 37),495 => (21, 37),496 => (22, 37),497 => (23, 37),498 => (24, 37),499 => (25, 37),500 => (26, 37),501 => (27, 37),502 => (34, 37),503 => (35, 37),504 => (41, 37),505 => (42, 37),506 => (46, 37),507 => (47, 37),508 => (48, 37),509 => (49, 37),510 => (50, 37),511 => (60, 37),512 => (61, 37),513 => (21, 38),514 => (22, 38),515 => (23, 38),516 => (24, 38),517 => (25, 38),518 => (26, 38),519 => (34, 38),520 => (35, 38),521 => (41, 38),522 => (42, 38),523 => (47, 38),524 => (48, 38),525 => (49, 38),526 => (50, 38),527 => (60, 38),528 => (61, 38),529 => (21, 39),530 => (22, 39),531 => (25, 39),532 => (26, 39),533 => (31, 39),534 => (32, 39),535 => (33, 39),536 => (34, 39),537 => (35, 39),538 => (36, 39),539 => (37, 39),540 => (38, 39),541 => (41, 39),542 => (42, 39),543 => (48, 39),544 => (49, 39),545 => (50, 39),546 => (52, 39),547 => (53, 39),548 => (54, 39),549 => (55, 39),550 => (56, 39),551 => (57, 39),552 => (58, 39),553 => (59, 39),554 => (60, 39),555 => (61, 39),556 => (21, 40),557 => (22, 40),558 => (25, 40),559 => (26, 40),560 => (31, 40),561 => (32, 40),562 => (33, 40),563 => (34, 40),564 => (35, 40),565 => (36, 40),566 => (37, 40),567 => (38, 40),568 => (41, 40),569 => (42, 40),570 => (49, 40),571 => (50, 40),572 => (52, 40),573 => (53, 40),574 => (54, 40),575 => (55, 40),576 => (56, 40),577 => (57, 40),578 => (58, 40),579 => (59, 40),580 => (60, 40),581 => (61, 40),others => (-1,-1));
constant player2WinsImage : coordinate_array (0 to FIXED_SCREEN_ELEMENTS - 1, 0 to 1) := (0 => (3, 19),1 => (4, 19),2 => (5, 19),3 => (6, 19),4 => (7, 19),5 => (8, 19),6 => (9, 19),7 => (10, 19),8 => (11, 19),9 => (12, 19),10 => (14, 19),11 => (15, 19),12 => (25, 19),13 => (26, 19),14 => (27, 19),15 => (28, 19),16 => (29, 19),17 => (30, 19),18 => (31, 19),19 => (32, 19),20 => (33, 19),21 => (34, 19),22 => (36, 19),23 => (37, 19),24 => (44, 19),25 => (45, 19),26 => (47, 19),27 => (48, 19),28 => (49, 19),29 => (50, 19),30 => (51, 19),31 => (52, 19),32 => (53, 19),33 => (54, 19),34 => (55, 19),35 => (56, 19),36 => (58, 19),37 => (59, 19),38 => (60, 19),39 => (61, 19),40 => (62, 19),41 => (63, 19),42 => (64, 19),43 => (65, 19),44 => (66, 19),45 => (67, 19),46 => (70, 19),47 => (71, 19),48 => (72, 19),49 => (73, 19),50 => (74, 19),51 => (75, 19),52 => (76, 19),53 => (3, 20),54 => (4, 20),55 => (5, 20),56 => (6, 20),57 => (7, 20),58 => (8, 20),59 => (9, 20),60 => (10, 20),61 => (11, 20),62 => (12, 20),63 => (14, 20),64 => (15, 20),65 => (25, 20),66 => (26, 20),67 => (27, 20),68 => (28, 20),69 => (29, 20),70 => (30, 20),71 => (31, 20),72 => (32, 20),73 => (33, 20),74 => (34, 20),75 => (36, 20),76 => (37, 20),77 => (38, 20),78 => (43, 20),79 => (44, 20),80 => (45, 20),81 => (47, 20),82 => (48, 20),83 => (49, 20),84 => (50, 20),85 => (51, 20),86 => (52, 20),87 => (53, 20),88 => (54, 20),89 => (55, 20),90 => (56, 20),91 => (58, 20),92 => (59, 20),93 => (60, 20),94 => (61, 20),95 => (62, 20),96 => (63, 20),97 => (64, 20),98 => (65, 20),99 => (66, 20),100 => (67, 20),101 => (69, 20),102 => (70, 20),103 => (71, 20),104 => (72, 20),105 => (73, 20),106 => (74, 20),107 => (75, 20),108 => (76, 20),109 => (77, 20),110 => (3, 21),111 => (4, 21),112 => (11, 21),113 => (12, 21),114 => (14, 21),115 => (15, 21),116 => (25, 21),117 => (26, 21),118 => (33, 21),119 => (34, 21),120 => (37, 21),121 => (38, 21),122 => (39, 21),123 => (42, 21),124 => (43, 21),125 => (44, 21),126 => (47, 21),127 => (48, 21),128 => (58, 21),129 => (59, 21),130 => (66, 21),131 => (67, 21),132 => (69, 21),133 => (70, 21),134 => (71, 21),135 => (75, 21),136 => (76, 21),137 => (77, 21),138 => (78, 21),139 => (3, 22),140 => (4, 22),141 => (11, 22),142 => (12, 22),143 => (14, 22),144 => (15, 22),145 => (25, 22),146 => (26, 22),147 => (33, 22),148 => (34, 22),149 => (38, 22),150 => (39, 22),151 => (40, 22),152 => (41, 22),153 => (42, 22),154 => (43, 22),155 => (47, 22),156 => (48, 22),157 => (58, 22),158 => (59, 22),159 => (66, 22),160 => (67, 22),161 => (75, 22),162 => (76, 22),163 => (77, 22),164 => (3, 23),165 => (4, 23),166 => (5, 23),167 => (6, 23),168 => (7, 23),169 => (8, 23),170 => (9, 23),171 => (10, 23),172 => (11, 23),173 => (12, 23),174 => (14, 23),175 => (15, 23),176 => (25, 23),177 => (26, 23),178 => (33, 23),179 => (34, 23),180 => (39, 23),181 => (40, 23),182 => (41, 23),183 => (42, 23),184 => (47, 23),185 => (48, 23),186 => (49, 23),187 => (50, 23),188 => (51, 23),189 => (52, 23),190 => (58, 23),191 => (59, 23),192 => (60, 23),193 => (61, 23),194 => (62, 23),195 => (63, 23),196 => (64, 23),197 => (65, 23),198 => (66, 23),199 => (67, 23),200 => (74, 23),201 => (75, 23),202 => (76, 23),203 => (3, 24),204 => (4, 24),205 => (5, 24),206 => (6, 24),207 => (7, 24),208 => (8, 24),209 => (9, 24),210 => (10, 24),211 => (11, 24),212 => (12, 24),213 => (14, 24),214 => (15, 24),215 => (25, 24),216 => (26, 24),217 => (27, 24),218 => (28, 24),219 => (29, 24),220 => (30, 24),221 => (31, 24),222 => (32, 24),223 => (33, 24),224 => (34, 24),225 => (40, 24),226 => (41, 24),227 => (47, 24),228 => (48, 24),229 => (49, 24),230 => (50, 24),231 => (51, 24),232 => (52, 24),233 => (58, 24),234 => (59, 24),235 => (60, 24),236 => (61, 24),237 => (62, 24),238 => (63, 24),239 => (64, 24),240 => (65, 24),241 => (66, 24),242 => (73, 24),243 => (74, 24),244 => (75, 24),245 => (3, 25),246 => (4, 25),247 => (14, 25),248 => (15, 25),249 => (25, 25),250 => (26, 25),251 => (27, 25),252 => (28, 25),253 => (29, 25),254 => (30, 25),255 => (31, 25),256 => (32, 25),257 => (33, 25),258 => (34, 25),259 => (40, 25),260 => (41, 25),261 => (47, 25),262 => (48, 25),263 => (58, 25),264 => (59, 25),265 => (63, 25),266 => (64, 25),267 => (65, 25),268 => (72, 25),269 => (73, 25),270 => (74, 25),271 => (3, 26),272 => (4, 26),273 => (14, 26),274 => (15, 26),275 => (25, 26),276 => (26, 26),277 => (33, 26),278 => (34, 26),279 => (40, 26),280 => (41, 26),281 => (47, 26),282 => (48, 26),283 => (58, 26),284 => (59, 26),285 => (64, 26),286 => (65, 26),287 => (66, 26),288 => (71, 26),289 => (72, 26),290 => (73, 26),291 => (3, 27),292 => (4, 27),293 => (14, 27),294 => (15, 27),295 => (16, 27),296 => (17, 27),297 => (18, 27),298 => (19, 27),299 => (20, 27),300 => (21, 27),301 => (22, 27),302 => (25, 27),303 => (26, 27),304 => (33, 27),305 => (34, 27),306 => (40, 27),307 => (41, 27),308 => (47, 27),309 => (48, 27),310 => (49, 27),311 => (50, 27),312 => (51, 27),313 => (52, 27),314 => (53, 27),315 => (54, 27),316 => (55, 27),317 => (56, 27),318 => (58, 27),319 => (59, 27),320 => (65, 27),321 => (66, 27),322 => (67, 27),323 => (70, 27),324 => (71, 27),325 => (72, 27),326 => (73, 27),327 => (74, 27),328 => (75, 27),329 => (76, 27),330 => (77, 27),331 => (78, 27),332 => (3, 28),333 => (4, 28),334 => (14, 28),335 => (15, 28),336 => (16, 28),337 => (17, 28),338 => (18, 28),339 => (19, 28),340 => (20, 28),341 => (21, 28),342 => (22, 28),343 => (25, 28),344 => (26, 28),345 => (33, 28),346 => (34, 28),347 => (40, 28),348 => (41, 28),349 => (47, 28),350 => (48, 28),351 => (49, 28),352 => (50, 28),353 => (51, 28),354 => (52, 28),355 => (53, 28),356 => (54, 28),357 => (55, 28),358 => (56, 28),359 => (58, 28),360 => (59, 28),361 => (66, 28),362 => (67, 28),363 => (69, 28),364 => (70, 28),365 => (71, 28),366 => (72, 28),367 => (73, 28),368 => (74, 28),369 => (75, 28),370 => (76, 28),371 => (77, 28),372 => (78, 28),373 => (19, 31),374 => (20, 31),375 => (27, 31),376 => (28, 31),377 => (31, 31),378 => (32, 31),379 => (33, 31),380 => (34, 31),381 => (35, 31),382 => (36, 31),383 => (37, 31),384 => (38, 31),385 => (41, 31),386 => (42, 31),387 => (49, 31),388 => (50, 31),389 => (52, 31),390 => (53, 31),391 => (54, 31),392 => (55, 31),393 => (56, 31),394 => (57, 31),395 => (58, 31),396 => (59, 31),397 => (60, 31),398 => (61, 31),399 => (19, 32),400 => (20, 32),401 => (27, 32),402 => (28, 32),403 => (31, 32),404 => (32, 32),405 => (33, 32),406 => (34, 32),407 => (35, 32),408 => (36, 32),409 => (37, 32),410 => (38, 32),411 => (41, 32),412 => (42, 32),413 => (43, 32),414 => (49, 32),415 => (50, 32),416 => (52, 32),417 => (53, 32),418 => (54, 32),419 => (55, 32),420 => (56, 32),421 => (57, 32),422 => (58, 32),423 => (59, 32),424 => (60, 32),425 => (61, 32),426 => (19, 33),427 => (20, 33),428 => (27, 33),429 => (28, 33),430 => (34, 33),431 => (35, 33),432 => (41, 33),433 => (42, 33),434 => (43, 33),435 => (44, 33),436 => (49, 33),437 => (50, 33),438 => (52, 33),439 => (53, 33),440 => (19, 34),441 => (20, 34),442 => (21, 34),443 => (23, 34),444 => (24, 34),445 => (26, 34),446 => (27, 34),447 => (28, 34),448 => (34, 34),449 => (35, 34),450 => (41, 34),451 => (42, 34),452 => (43, 34),453 => (44, 34),454 => (45, 34),455 => (49, 34),456 => (50, 34),457 => (52, 34),458 => (53, 34),459 => (20, 35),460 => (21, 35),461 => (23, 35),462 => (24, 35),463 => (26, 35),464 => (27, 35),465 => (34, 35),466 => (35, 35),467 => (41, 35),468 => (42, 35),469 => (44, 35),470 => (45, 35),471 => (46, 35),472 => (49, 35),473 => (50, 35),474 => (52, 35),475 => (53, 35),476 => (54, 35),477 => (55, 35),478 => (56, 35),479 => (57, 35),480 => (58, 35),481 => (59, 35),482 => (60, 35),483 => (61, 35),484 => (20, 36),485 => (21, 36),486 => (22, 36),487 => (23, 36),488 => (24, 36),489 => (25, 36),490 => (26, 36),491 => (27, 36),492 => (34, 36),493 => (35, 36),494 => (41, 36),495 => (42, 36),496 => (45, 36),497 => (46, 36),498 => (47, 36),499 => (49, 36),500 => (50, 36),501 => (52, 36),502 => (53, 36),503 => (54, 36),504 => (55, 36),505 => (56, 36),506 => (57, 36),507 => (58, 36),508 => (59, 36),509 => (60, 36),510 => (61, 36),511 => (20, 37),512 => (21, 37),513 => (22, 37),514 => (23, 37),515 => (24, 37),516 => (25, 37),517 => (26, 37),518 => (27, 37),519 => (34, 37),520 => (35, 37),521 => (41, 37),522 => (42, 37),523 => (46, 37),524 => (47, 37),525 => (48, 37),526 => (49, 37),527 => (50, 37),528 => (60, 37),529 => (61, 37),530 => (21, 38),531 => (22, 38),532 => (23, 38),533 => (24, 38),534 => (25, 38),535 => (26, 38),536 => (34, 38),537 => (35, 38),538 => (41, 38),539 => (42, 38),540 => (47, 38),541 => (48, 38),542 => (49, 38),543 => (50, 38),544 => (60, 38),545 => (61, 38),546 => (21, 39),547 => (22, 39),548 => (25, 39),549 => (26, 39),550 => (31, 39),551 => (32, 39),552 => (33, 39),553 => (34, 39),554 => (35, 39),555 => (36, 39),556 => (37, 39),557 => (38, 39),558 => (41, 39),559 => (42, 39),560 => (48, 39),561 => (49, 39),562 => (50, 39),563 => (52, 39),564 => (53, 39),565 => (54, 39),566 => (55, 39),567 => (56, 39),568 => (57, 39),569 => (58, 39),570 => (59, 39),571 => (60, 39),572 => (61, 39),573 => (21, 40),574 => (22, 40),575 => (25, 40),576 => (26, 40),577 => (31, 40),578 => (32, 40),579 => (33, 40),580 => (34, 40),581 => (35, 40),582 => (36, 40),583 => (37, 40),584 => (38, 40),585 => (41, 40),586 => (42, 40),587 => (49, 40),588 => (50, 40),589 => (52, 40),590 => (53, 40),591 => (54, 40),592 => (55, 40),593 => (56, 40),594 => (57, 40),595 => (58, 40),596 => (59, 40),597 => (60, 40),598 => (61, 40), others => (-1,-1));

begin 

process(clk)

variable hMatrix, vMatrix : integer := 0;
variable draw : std_logic := '0';

variable is_element : std_logic := '0';
variable is_special : std_logic := '0';
variable is_player1 : std_logic := '0';
variable is_player2 : std_logic := '0';

begin

	if(rising_edge(clk)) then
		if(draw = '1') then
			if(gameStarted = '0') then
				hMatrix := (hpos - H_OFFSET)/PIXEL_SIZE;
				vMatrix := (vpos - V_OFFSET)/PIXEL_SIZE;
				if((hpos - H_OFFSET) MOD PIXEL_SIZE = 0 or (vpos - V_OFFSET) MOD PIXEL_SIZE = 0) then
					r <= (others => '0');
					g <= (others => '0');
					b <= (others => '0');
				else
					is_element := '0';
					for i in 0 to FIXED_SCREEN_ELEMENTS - 1 loop
						if(vMatrix = gameStartImage(i, 1)) then
							if(hMatrix = gameStartImage(i,0)) then
								is_element := '1';
							end if;
						end if;
					end loop;
					
					if(is_element = '1') then
						r <= (others => '1');
						g <= (others => '1');
						b <= (others => '1');
					else
						r <= (0 => '1', others => '0');
						g <= (0 => '1', others => '0');
						b <= (0 => '1', others => '0');
					end if;
				end if;
			elsif(player1won = '1') then
				hMatrix := (hpos - H_OFFSET)/PIXEL_SIZE;
				vMatrix := (vpos - V_OFFSET)/PIXEL_SIZE;
				if((hpos - H_OFFSET) REM PIXEL_SIZE = 0 or (vpos - V_OFFSET) REM PIXEL_SIZE = 0) then
					r <= (others => '0');
					g <= (others => '0');
					b <= (others => '0');
				else
					is_element := '0';
					for i in 0 to FIXED_SCREEN_ELEMENTS - 1 loop
						if(vMatrix = player1winsImage(i, 1)) then
							if(hMatrix = player1winsImage(i,0)) then
								is_element := '1';
							end if;
						end if;
						if(is_element = '1') then
							r <= (others => '1');
							g <= (others => '1');
							b <= (others => '1');
						else
							r <= (0 => '1', others => '0');
							g <= (0 => '1', others => '0');
							b <= (0 => '1', others => '0');
						end if;
					end loop;
				end if;
			elsif(player2won = '1') then
				hMatrix := (hpos - H_OFFSET)/PIXEL_SIZE;
				vMatrix := (vpos - V_OFFSET)/PIXEL_SIZE;
				if((hpos - H_OFFSET) REM PIXEL_SIZE = 0 or (vpos - V_OFFSET) REM PIXEL_SIZE = 0) then
					r <= (others => '0');
					g <= (others => '0');
					b <= (others => '0');
				else
					is_element := '0';
					for i in 0 to FIXED_SCREEN_ELEMENTS - 1 loop
						if(vMatrix = player2winsImage(i, 1)) then
							if(hMatrix = player2winsImage(i,0)) then
								is_element := '1';
							end if;
						end if;						
						if(is_element = '1') then
							r <= (others => '1');
							g <= (others => '1');
							b <= (others => '1');
						else
							r <= (0 => '1', others => '0');
							g <= (0 => '1', others => '0');
							b <= (0 => '1', others => '0');
						end if;
					end loop;
				end if;
			elsif(gameStarted = '1' and player1won = '0' and player2won = '0') then
				hMatrix := (hpos - H_OFFSET)/PIXEL_SIZE;
				vMatrix := (vpos - V_OFFSET)/PIXEL_SIZE;
				if((hpos - H_OFFSET) REM PIXEL_SIZE = 0 or (vpos - V_OFFSET) REM PIXEL_SIZE = 0) then
					r <= (others => '0');
					g <= (others => '0');
					b <= (others => '0');
				else
					is_player1 := '0';
					for i in 0 to MAX_ELEMENTS - 1 loop
						if(vMatrix = player1(i, 1)) then
							if(hMatrix = player1(i,0)) then
								if(circleImage((hpos - H_OFFSET) REM PIXEL_SIZE, (vpos - V_OFFSET) REM PIXEL_SIZE) = '0') then
									is_player1 := '1';
								end if;
							end if;
						end if;
					end loop;	
					is_player2 := '0';
					for i in 0 to MAX_ELEMENTS - 1 loop
						if(vMatrix = player2(i, 1)) then
							if(hMatrix = player2(i,0)) then
								if(circleImage((hpos - H_OFFSET) REM PIXEL_SIZE, (vpos - V_OFFSET) REM PIXEL_SIZE) = '0') then
									is_player2 := '1';
								end if;
							end if;
						end if;
					end loop;
							
					is_element := '0';
					if(vMatrix = apple_position(1)) then
						if(hMatrix = apple_position(0)) then
							if(circleImage((hpos - H_OFFSET) REM PIXEL_SIZE, (vpos - V_OFFSET) REM PIXEL_SIZE) = '0') then	
								is_element := '1';
							end if;
						end if;
					end if;
					is_special := '0';
					if(vMatrix = special_position(1)) then
						if(hMatrix = special_position(0)) then
							if(circleImage((hpos - H_OFFSET) REM PIXEL_SIZE, (vpos - V_OFFSET) REM PIXEL_SIZE) = '0') then	
								is_special := '1';
							end if;
						end if;
					end if;
					
					if(is_player1 = '1') then
						r <= (others => '1');
						g <= (others => '0');
						b <= (others => '1');
					elsif(is_player2 = '1') then
						r <= (others => '0');
						g <= (others => '0');
						b <= (others => '1');
					elsif(is_special = '1') then
						r <= (others => '0');
						g <= (others => '1');
						b <= (others => '0');
					elsif(is_element = '1') then
						r <= (others => '1');
						g <= (others => '1');
						b <= (others => '1');
					else
						r <= (0 => '1', others => '0');
						g <= (0 => '1', others => '0');
						b <= (0 => '1', others => '0');
					end if;
				end if;
			end if;
		else	
				r <= (0 => '1',others => '0');
				g <= (0 => '1',others => '0');
				b <= (0 => '1',others => '0');
		end if;
		if(hpos < H_OFFSET + H_SIZE) then
			hpos<= hpos +1;
		else
			hpos<= 0;
			if(vpos < 1066) then
				vpos<= vpos + 1;
			else
				vpos <= 0;
			end if;
		end if;
	end if;
	if(hpos >H_FP and hpos <H_FP + H_SYNCP) then
		hsync <= '0';
	else
		hsync <= '1';
	end if;
	if(vpos > 0 and vpos < V_FP + V_SYNCP) then
		vsync <= '0';
	else
		vsync <= '1';
	end if;
	if((hpos > 0 and hpos < H_OFFSET) or (vpos >0 and vpos <V_OFFSET)) then
		r<= (others => '0');
		g<= (others => '0');
		b<= (others => '0');
		draw := '0';
	else
		draw := '1';
	end if;
end process;

end architecture;